(a+bi)*(c+di)=(ac-bd)+(ad+bc)i
4 multiplys, 3 adds

optimization:
A = (a+b)*c
B = (c+d)*b
C = (b-a)*d
(a+bi)*(c+di) = (A-B)+(B-C)i
3 multiplys, 6 adds
Add is much faster than multiply.
